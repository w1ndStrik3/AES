library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package heap_arr_pkg is
    type round_key_t is array(0 to 14) of std_logic_vector(127 downto 0);
end; 